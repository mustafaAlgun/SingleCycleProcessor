library verilog;
use verilog.vl_types.all;
entity SingleCycleProcessor_tb is
end SingleCycleProcessor_tb;
